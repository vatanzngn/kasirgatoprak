// Onbellek ile alakalı yapilandirma
`include "sentez_tanimlari.vh"

`define BOLME_HER_CEVRIM_BIT_SAYISI 1
`define ONBELLEK_SATIR_SOZCUK_SAYISI 4
`define L1_BUYRUK_ONBELLEK_YOL_SAYISI 2
`define L1_BUYRUK_ONBELLEK_YOL_SATIR_SAYISI 128
`define L1_VERI_ONBELLEK_YOL_SAYISI 2
`define L1_VERI_ONBELLEK_YOL_SATIR_SAYISI 128
`define ADRES_ONEMSIZ_BIT_SAYISI 2
`define BASLANGIC_ADRESI 32'h8000_0000
`define BITIS_ADRESI 32'h8100_0000
`define YENI_RAM_MODELI_GECIKME 0
`define RAM_SATIR_SAYISI 512
`define RAM_SATIR_SOZCUK_SAYISI 4
`define WB_SLAVE_SAYISI 1

//`define WB_UART
