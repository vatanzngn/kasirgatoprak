package oncoz_pkg;

   typedef enum logic [1:0] {
      DALLANMA,
      JAL,
      JALR,
      DALLANMA_YOK
   } dallanma_turu_t;

endpackage : oncoz_pkg
