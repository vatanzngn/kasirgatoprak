`define USE_SRAM
`define BASYS3
//`define NEXYS7
//`define VCU108
`define SPIKE_DIFF
`define FPU // FPUyu acar
`define DEBUG
//`define REM_IP // ipleri kaldırır
//`define YUKSEK_BOYUT_UART_FIFO

