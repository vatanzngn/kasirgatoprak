`define NOP 32'h00000013

`define SOZCUK_GENISLIGI_BIT 32
`define ADRES_GENISLIGI_BIT 32

`define BELLEK_KONTROL_SINYALI_BIT 9
`define MASKE_GENISLIGI_BIT 4

`define HIGH 1
`define LOW 0

// CSR_SABITLERI
`define CSR_MOD_BITIS 11
`define CSR_MOD_BASLANGIC 10

`define CSR_DUZEY_BASLANGIC 8
`define CSR_DUZEY_BITIS 9

`define CSR_DUZEY_UNPRIV 2'b00
`define CSR_DUZEY_SUPERV 2'b01
`define CSR_DUZEY_HYPERV 2'b10
`define CSR_DUZEY_MACHINE 2'b11

`define CSR_MOD_SALT_OKUNUR 2'b11
`define CSR_MOD_YAZILABILIR 2'b00 || 2'b01 || 2'b10

`define CSR_WR_WPRI 2'b00 // YAZMAYA VE OKUMAYA IZIN VER YAZILIM OKUNAN VERIYI UMURSAMAMALI
`define CSR_WR_WLRL 2'b01 // YAZARKEN VE OKURKEN VERILEN GIRDI GECERLI OLMASI ZORUNLU ILLEGAL INSTRUCTION FIRLATILABILIR AMA ZORUNLU DEGIL
`define CSR_WR_WARL 2'b1x // YAZMAYA IZIN VERMIŞ GİBİ GOSTER AMA SADECE LEGAL DEGER OKUNABILIR

// MACHINE_MODE Denetim Durum Yazmaç adresleri
`define CSR_ADDR_MSTATUS 12'h300
`define CSR_ADDR_MISA 12'h301
`define CSR_ADDR_MEDELEG 12'h302
`define CSR_ADDR_MIDELEG 12'h303
`define CSR_ADDR_MIE 12'h304
`define CSR_ADDR_MTVEC 12'h305
`define CSR_ADDR_MCOUNTEREN 12'h306
`define CSR_ADDR_MSTATUSH 12'h310
`define CSR_ADDR_MSCRATCH 12'h340
`define CSR_ADDR_MEPC 12'h341
`define CSR_ADDR_MCAUSE 12'h342
`define CSR_ADDR_MTVAL 12'h343
`define CSR_ADDR_MIP 12'h344
`define CSR_ADDR_MTINST 12'h34A
`define CSR_ADDR_MTVAL2 12'h34B
`define CSR_ADDR_MCYCLE 12'hB00
`define CSR_ADDR_MINSTRET 12'hB02
`define CSR_ADDR_MVENVCFG 12'h30A
`define CSR_ADDR_MVENVCFGH 12'h31A
`define CSR_ADDR_MHPMCOUNTER3 12'hB03
`define CSR_ADDR_MHPMCOUNTER4 12'hB04
`define CSR_ADDR_MHPMCOUNTER5 12'hB05
`define CSR_ADDR_MHPMCOUNTER6 12'hB06
`define CSR_ADDR_MHPMCOUNTER7 12'hB07
`define CSR_ADDR_MHPMCOUNTER8 12'hB08
`define CSR_ADDR_MHPMCOUNTER9 12'hB09
`define CSR_ADDR_MHPMCOUNTER10 12'hB0A
`define CSR_ADDR_MHPMCOUNTER11 12'hB0B
`define CSR_ADDR_MHPMCOUNTER12 12'hB0C
`define CSR_ADDR_MHPMCOUNTER13 12'hB0D
`define CSR_ADDR_MHPMCOUNTER14 12'hB0E
`define CSR_ADDR_MHPMCOUNTER15 12'hB0F
`define CSR_ADDR_MHPMCOUNTER16 12'hB10
`define CSR_ADDR_MHPMCOUNTER17 12'hB11
`define CSR_ADDR_MHPMCOUNTER18 12'hB12
`define CSR_ADDR_MHPMCOUNTER19 12'hB13
`define CSR_ADDR_MHPMCOUNTER20 12'hB14
`define CSR_ADDR_MHPMCOUNTER21 12'hB15
`define CSR_ADDR_MHPMCOUNTER22 12'hB16
`define CSR_ADDR_MHPMCOUNTER23 12'hB17
`define CSR_ADDR_MHPMCOUNTER24 12'hB18
`define CSR_ADDR_MHPMCOUNTER25 12'hB19
`define CSR_ADDR_MHPMCOUNTER26 12'hB1A
`define CSR_ADDR_MHPMCOUNTER27 12'hB1B
`define CSR_ADDR_MHPMCOUNTER28 12'hB1C
`define CSR_ADDR_MHPMCOUNTER29 12'hB1D
`define CSR_ADDR_MHPMCOUNTER30 12'hB1E
`define CSR_ADDR_MHPMCOUNTER31 12'hB1F
`define CSR_ADDR_MCOUNTINHIBIT 12'h320
`define CSR_ADDR_MHPEVENT3 12'h323
`define CSR_ADDR_MHPEVENT4 12'h324
`define CSR_ADDR_MHPEVENT5 12'h325
`define CSR_ADDR_MHPEVENT6 12'h326
`define CSR_ADDR_MHPEVENT7 12'h327
`define CSR_ADDR_MHPEVENT8 12'h328
`define CSR_ADDR_MHPEVENT9 12'h329
`define CSR_ADDR_MHPEVENT10 12'h32A
`define CSR_ADDR_MHPEVENT11 12'h32B
`define CSR_ADDR_MHPEVENT12 12'h32C
`define CSR_ADDR_MHPEVENT13 12'h32D
`define CSR_ADDR_MHPEVENT14 12'h32E
`define CSR_ADDR_MHPEVENT15 12'h32F
`define CSR_ADDR_MHPEVENT16 12'h330
`define CSR_ADDR_MHPEVENT17 12'h331
`define CSR_ADDR_MHPEVENT18 12'h332
`define CSR_ADDR_MHPEVENT19 12'h333
`define CSR_ADDR_MHPEVENT20 12'h334
`define CSR_ADDR_MHPEVENT21 12'h335
`define CSR_ADDR_MHPEVENT22 12'h336
`define CSR_ADDR_MHPEVENT23 12'h337
`define CSR_ADDR_MHPEVENT24 12'h338
`define CSR_ADDR_MHPEVENT25 12'h339
`define CSR_ADDR_MHPEVENT26 12'h33A
`define CSR_ADDR_MHPEVENT27 12'h33B
`define CSR_ADDR_MHPEVENT28 12'h33C
`define CSR_ADDR_MHPEVENT29 12'h33D
`define CSR_ADDR_MHPEVENT30 12'h33E
`define CSR_ADDR_MHPEVENT31 12'h33F
`define CSR_ADDR_MCYCLEH 12'hB80
`define CSR_ADDR_MINSTRETH 12'hB82
`define CSR_ADDR_MHPMCOUNTER3H 12'hB83
`define CSR_ADDR_MHPMCOUNTER4H 12'hB84
`define CSR_ADDR_MHPMCOUNTER5H 12'hB85
`define CSR_ADDR_MHPMCOUNTER6H 12'hB86
`define CSR_ADDR_MHPMCOUNTER7H 12'hB87
`define CSR_ADDR_MHPMCOUNTER8H 12'hB88
`define CSR_ADDR_MHPMCOUNTER9H 12'hB89
`define CSR_ADDR_MHPMCOUNTER10H 12'hB8A
`define CSR_ADDR_MHPMCOUNTER11H 12'hB8B
`define CSR_ADDR_MHPMCOUNTER12H 12'hB8C
`define CSR_ADDR_MHPMCOUNTER13H 12'hB8D
`define CSR_ADDR_MHPMCOUNTER14H 12'hB8E
`define CSR_ADDR_MHPMCOUNTER15H 12'hB8F
`define CSR_ADDR_MHPMCOUNTER16H 12'hB90
`define CSR_ADDR_MHPMCOUNTER17H 12'hB91
`define CSR_ADDR_MHPMCOUNTER18H 12'hB92
`define CSR_ADDR_MHPMCOUNTER19H 12'hB93
`define CSR_ADDR_MHPMCOUNTER20H 12'hB94
`define CSR_ADDR_MHPMCOUNTER21H 12'hB95
`define CSR_ADDR_MHPMCOUNTER22H 12'hB96
`define CSR_ADDR_MHPMCOUNTER23H 12'hB97
`define CSR_ADDR_MHPMCOUNTER24H 12'hB98
`define CSR_ADDR_MHPMCOUNTER25H 12'hB99
`define CSR_ADDR_MHPMCOUNTER26H 12'hB9A
`define CSR_ADDR_MHPMCOUNTER27H 12'hB9B
`define CSR_ADDR_MHPMCOUNTER28H 12'hB9C
`define CSR_ADDR_MHPMCOUNTER29H 12'hB9D
`define CSR_ADDR_MHPMCOUNTER30H 12'hB9E
`define CSR_ADDR_MHPMCOUNTER31H 12'hB9F
`define CSR_ADDR_MVENDORID 12'hF11
`define CSR_ADDR_MARCHID 12'hF12
`define CSR_ADDR_MIMPID 12'hF13
`define CSR_ADDR_MHARTID 12'hF14
`define CSR_ADDR_MCONFIGPTR 12'hF15
`define CSR_ADDR_PMPCFG0 12'h3A0
`define CSR_ADDR_PMPCFG1 12'h3A1
`define CSR_ADDR_PMPCFG2 12'h3A2
`define CSR_ADDR_PMPCFG3 12'h3A3
`define CSR_ADDR_PMPADDR0 12'h3B0
`define CSR_ADDR_PMPADDR1 12'h3B1
`define CSR_ADDR_PMPADDR2 12'h3B2
`define CSR_ADDR_PMPADDR3 12'h3B3
`define CSR_ADDR_PMPADDR4 12'h3B4
`define CSR_ADDR_PMPADDR5 12'h3B5
`define CSR_ADDR_PMPADDR6 12'h3B6
`define CSR_ADDR_PMPADDR7 12'h3B7
`define CSR_ADDR_PMPADDR8 12'h3B8
`define CSR_ADDR_PMPADDR9 12'h3B9
`define CSR_ADDR_PMPADDR10 12'h3BA
`define CSR_ADDR_PMPADDR11 12'h3BB
`define CSR_ADDR_PMPADDR12 12'h3BC
`define CSR_ADDR_PMPADDR13 12'h3BD
`define CSR_ADDR_PMPADDR14 12'h3BE
`define CSR_ADDR_PMPADDR15 12'h3BF

//USER_MODE uygulanacak CSR'lar FP-CSRs, C00-C02 (cycle, time, instrent)
//FPU ile ilgili alan
`define CSR_FPU_BASLANGIC 12'h001
`define CSR_FPU_BITIS 12'h001

`define CSR_ADDR_FFLAGS 12'h001
`define CSR_ADDR_FRM 12'h002
`define CSR_ADDR_FCSR 12'h003

`define CSR_ADDR_FFLAGS_H 12'h004

//USER MODE IMPLEMENT EDILEN CSRLAR
`define CSR_ADDR_CYCLE 12'hC00
`define CSR_ADDR_TIME 12'hC01
`define CSR_ADDR_INSTRET 12'hC02
`define CSR_ADDR_CYCLEH 12'hC80
`define CSR_ADDR_TIMEH 12'hC81
`define CSR_ADDR_INSTRETH 12'hC82
`define CSR_ADDR_HPMCOUNTER3 12'hC03
`define CSR_ADDR_HPMCOUNTER4 12'hC04
`define CSR_ADDR_HPMCOUNTER5 12'hC05
`define CSR_ADDR_HPMCOUNTER6 12'hC06

`define CSR_ADDR_HPMCOUNTER3H 12'hC83
`define CSR_ADDR_HPMCOUNTER4H 12'hC84
`define CSR_ADDR_HPMCOUNTER5H 12'hC85
`define CSR_ADDR_HPMCOUNTER6H 12'hC86
//DEBUG MODE IMPLEMENT EDILEN CSRLAR
`define CSR_ADDR_DCSR 12'h7B0
`define CSR_ADDR_DPC 12'h7B1
`define CSR_ADDR_DSCRATCH0 12'h7B2
`define CSR_ADDR_DSCRATCH1 12'h7B3

`define CSR_FUNCT3_CSRRW 3'b001
`define CSR_FUNCT3_CSRRS 3'b010
`define CSR_FUNCT3_CSRRC 3'b011
`define CSR_FUNCT3_CSRRWI 3'b101
`define CSR_FUNCT3_CSRRSI 3'b110
`define CSR_FUNCT3_CSRRCI 3'b111

`define CSR_MRET_FUNCT12 12'b001100000010
`define CSR_MRET_FUNCT3 3'b000

`define CSR_PRIV_BITIS 9
`define CSR_PRIV_BASLANGIC 8 
`define CSR_PRIV_USER 2'b00
`define CSR_PRIV_SV 2'b01
`define CSR_PRIV_HV 2'b10
`define CSR_PRIV_MACHINE 2'b11

`define MXL 1 // MXL değişince MXLEN guncellenmeli!!
`define MXL_MOD `CSR_MOD_SALT_OKUNUR

`define MXLEN 32 // MXL değişirse MXLEN güncellenmeli!!
`define CSR_MVENDOR_BIT 32
`define CSR_MVENDOR_DEGER 32'h0

`define CSR_MARCHID_BIT `MXLEN
`define CSR_MARCHID_DEGER 32'h0

`define CSR_MIMPID_BIT `MXLEN
`define CSR_MIMPID_DEGER 32'h001

`define CSR_MHARTID_BIT `MXLEN
`define CSR_MHARTID_DEGER 32'h0 // bir hartın 0 idli olması zorunlu, tek donanımsal threade sahip olduğumuzdan hardcoded 0

`define CSR_MCONFIGPTR_BIT `MXLEN
`define CSR_MCONFIGPTR_DEGER 32'h6000_0000 // umarım dolu degildir.

`define CSR_MSTATUS_BIT 32
`define CSR_MSTATUSH_BIT 32

`define CSR_MCYCLE_BIT 32
`define CSR_MCYCLEH_BIT 32

`define CSR_MISA_A 0
`define CSR_MISA_B 1
`define CSR_MISA_F 5
`define CSR_MISA_M 12

`define EXC_IAM 4'b0001
`define EXC_IAF 4'b0010
`define EXC_II 4'b0011
`define EXC_BP 4'b0100
`define EXC_LAM 4'b0101
`define EXC_LAF 4'b0110
`define EXC_SAM 4'b0111
`define EXC_SAF 4'b1000
`define EXC_ECALL 4'b1001
`define EXC_MRET 4'b1010

`define NOT_EXC_INV 4'b1111

`define EXC_IAM_CODE 0
`define EXC_IAF_CODE 1
`define EXC_II_CODE 2
`define EXC_BP_CODE 3
`define EXC_LAM_CODE 4
`define EXC_LAF_CODE 5
`define EXC_SAM_CODE 6
`define EXC_SAF_CODE 7
`define EXC_ECALL_CODE 11

`define MTVEC_MODE_DIRECT 0
`define MTVEC_MODE_VECTORED 1

////////////////////////////
`define CEVRE_BIRIM_BASLANGIC 32'h20_000_000
`define UART_BASLANGIC_ADRESI 32'h20_000_000
`define UART_BITIS_ADRESI 32'h20_000_00c

// gereksiz ama ek cevre birim baglanabilir diye birakiyorum
`define CEVRE_BIRIM_BITIS 32'h20_000_04c

`define UART_RX_FIFO_UZUNLUK 32
`define UART_TX_FIFO_UZUNLUK 32
`define UART_FIFO_GENISLIK 8
