// Kasırga - Toprak Buyruklar

// RV32I Buyrukları
`define I_LUI 32'b?????????????????????????0110111
`define I_AUIPC 32'b?????????????????????????0010111
`define I_JAL 32'b?????????????????????????1101111
`define I_JALR 32'b?????????????????000?????1100111
`define I_BEQ 32'b?????????????????000?????1100011
`define I_BNE 32'b?????????????????001?????1100011
`define I_BLT 32'b?????????????????100?????1100011
`define I_BGE 32'b?????????????????101?????1100011
`define I_BLTU 32'b?????????????????110?????1100011
`define I_BGEU 32'b?????????????????111?????1100011
`define I_LB 32'b?????????????????000?????0000011
`define I_LH 32'b?????????????????001?????0000011
`define I_LW 32'b?????????????????010?????0000011
`define I_LBU 32'b?????????????????100?????0000011
`define I_LHU 32'b?????????????????101?????0000011
`define I_SB 32'b?????????????????000?????0100011
`define I_SH 32'b?????????????????001?????0100011
`define I_SW 32'b?????????????????010?????0100011
`define I_ADDI 32'b?????????????????000?????0010011
`define I_SLTI 32'b?????????????????010?????0010011
`define I_SLTIU 32'b?????????????????011?????0010011
`define I_XORI 32'b?????????????????100?????0010011
`define I_ORI 32'b?????????????????110?????0010011
`define I_ANDI 32'b?????????????????111?????0010011
`define I_SLLI 32'b0000000??????????001?????0010011
`define I_SRLI 32'b0000000??????????101?????0010011
`define I_SRAI 32'b0100000??????????101?????0010011
`define I_ADD 32'b0000000??????????000?????0110011
`define I_SUB 32'b0100000??????????000?????0110011
`define I_SLL 32'b0000000??????????001?????0110011
`define I_SLT 32'b0000000??????????010?????0110011
`define I_SLTU 32'b0000000??????????011?????0110011
`define I_XOR 32'b0000000??????????100?????0110011
`define I_SRL 32'b0000000??????????101?????0110011
`define I_SRA 32'b0100000??????????101?????0110011
`define I_OR 32'b0000000??????????110?????0110011
`define I_AND 32'b0000000??????????111?????0110011
// RV32M Buyrukları//
`define I_MUL 32'b0000001??????????000?????0110011
`define I_MULH 32'b0000001??????????001?????0110011
`define I_MULHSU 32'b0000001??????????010?????0110011
`define I_MULHU 32'b0000001??????????011?????0110011
`define I_DIV 32'b0000001??????????100?????0110011
`define I_DIVU 32'b0000001??????????101?????0110011
`define I_REM 32'b0000001??????????110?????0110011
`define I_REMU 32'b0000001??????????111?????0110011
// RV32A Buyrukları//                                     
`define I_SC_W 32'b00011????????????010?????0101111
`define I_AMOSWAP_W 32'b00001????????????010?????0101111
`define I_AMOADD_W 32'b00000????????????010?????0101111
`define I_AMOXOR_W 32'b00100????????????010?????0101111
`define I_AMOAND_W 32'b01100????????????010?????0101111
`define I_AMOOR_W 32'b01000????????????010?????0101111
`define I_AMOMIN_W 32'b10000????????????010?????0101111
`define I_AMOMAX_W 32'b10100????????????010?????0101111
`define I_AMOMINU_W 32'b11000????????????010?????0101111
`define I_AMOMAXU_W 32'b11100????????????010?????0101111
//RV32F Buyrukları//
`define I_FLW 32'b?????????????????010?????0000111
`define I_FSW 32'b?????????????????010?????0100111
`define I_FMADD_S 32'b?????00??????????????????1000011
`define I_FMSUB_S 32'b?????00??????????????????1000111
`define I_FNMSUB_S 32'b?????00??????????????????1001011
`define I_FNMADD_S 32'b?????00??????????????????1001111
`define I_FADD_S 32'b0000000??????????????????1010011
`define I_FSUB_S 32'b0000100??????????????????1010011
`define I_FMUL_S 32'b0001000??????????????????1010011
`define I_FDIV_S 32'b0001100??????????????????1010011
`define I_FSQRT_S 32'b010110000000?????????????1010011
`define I_FSGNJ_S 32'b0010000??????????000?????1010011
`define I_FSGNJN_S 32'b0010000??????????001?????1010011
`define I_FSGNJX_S 32'b0010000??????????010?????1010011
`define I_FMIN_S 32'b0010100??????????000?????1010011
`define I_FMAX_S 32'b0010100??????????001?????1010011
`define I_FCVT_W_S 32'b110000000000?????????????1010011
`define I_FCVT_WU_S 32'b110000000001?????????????1010011
`define I_FMV_X_W 32'b111000000000?????000?????1010011
`define I_FEQ_S 32'b1010000??????????010?????1010011
`define I_FLT_S 32'b1010000??????????001?????1010011
`define I_FLE_S 32'b1010000??????????000?????1010011
`define I_FCLASS_S 32'b111000000000?????001?????1010011
`define I_FCVT_S_W 32'b110100000000?????????????1010011
`define I_FCVT_S_WU 32'b110100000001?????????????1010011
`define I_FMV_W_X 32'b111100000000?????000?????1010011
// RV32B Buyrukları
`define I_ADDN 32'b0100000??????????111?????0110011
`define I_CLMUL 32'b0000101??????????001?????0110011
`define I_CLMULH 32'b0000101??????????011?????0110011
`define I_CLMULR 32'b0000101??????????010?????0110011
`define I_CLZ 32'b011000000000?????001?????0010011 
`define I_CPOP 32'b011000000010?????001?????0010011
`define I_CTZ 32'b011000000001?????001?????0010011 
`define I_MAX 32'b0000101??????????110?????0110011
`define I_MAXU 32'b0000101??????????111?????0110011
`define I_MIN 32'b0000101??????????100?????0110011
`define I_MINU 32'b0000101??????????101?????0110011
`define I_ORC_B 32'b001010000111?????101?????0010011
`define I_ORN 32'b0100000??????????110?????0110011
`define I_REV8 32'b011010011000?????101?????0010011
`define I_ROL 32'b0110000??????????001?????0110011
`define I_ROR 32'b0110000??????????101?????0110011
`define I_RORI 32'b01100????????????101?????0010011
`define I_BCLR 32'b0100100??????????001?????0110011
`define I_BCLRI 32'b01001????????????001?????0010011
`define I_BEXT 32'b0100100??????????101?????0110011
`define I_BEXTI 32'b01001????????????101?????0010011
`define I_BINV 32'b0110100??????????001?????0110011
`define I_BINVI 32'b01101????????????001?????0010011
`define I_BSET 32'b0010100??????????001?????0110011
`define I_BSETI 32'b00101????????????001?????0010011
`define I_SEXT_B 32'b011000000100?????001?????0010011
`define I_SEXT_H 32'b011000000101?????001?????0010011
`define I_SH1ADD 32'b0010000??????????010?????0110011
`define I_SH2ADD 32'b0010000??????????100?????0110011
`define I_SH3ADD 32'b0010000??????????110?????0110011
`define I_XNOR 32'b0100000??????????100?????0110011
`define I_ZEXT_H 32'b000010000000?????100?????0110011

